package test_pkg; 

	import uvm_pkg::*;

	`include "uvm_macros.svh"

	`include "src_agent.sv"
	`include "dst_agent.sv"

	`include "env.sv"

	`include "test.sv"

endpackage

